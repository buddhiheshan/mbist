module controller #(
    parameters
) (
    ports
);
    
endmodule