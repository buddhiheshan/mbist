module decoder #(
    parameters
) (
    ports
);
    
endmodule