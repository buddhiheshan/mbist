module tb_bist ();
    
endmodule